`include "mips_defines.v"

`define ADDR_WIDTH 9
`define INSTR_WIDTH 32
`define NUM_INSTR 512

module irom(clk, addr, dout);
    input clk;
    input [`ADDR_WIDTH-1:0] addr;
    output reg [`INSTR_WIDTH-1:0] dout;
    
    wire [`INSTR_WIDTH-1:0] memory [`NUM_INSTR-1:0];
    
    always @(posedge clk)
        dout <= memory[addr];

assign memory[0] = {`SPECIAL, `ZERO, `ZERO, `SP, 5'd0, `ADD};
assign memory[1] = {`ADDI, `ZERO, `T0, 16'd39};
assign memory[2] = {`SW, `SP, `T0, 16'd0};
assign memory[3] = {`ADDI, `ZERO, `T0, 16'd29};
assign memory[4] = {`SW, `SP, `T0, 16'd4};
assign memory[5] = {`ADDI, `ZERO, `T0, 16'd0};
assign memory[6] = {`SW, `SP, `T0, 16'd8};
assign memory[7] = {`ADDI, `ZERO, `T0, 16'd2};
assign memory[8] = {`SW, `SP, `T0, 16'd12};
assign memory[9] = {`ADDI, `ZERO, `T0, 16'd4};
assign memory[10] = {`SW, `SP, `T0, 16'd16};
assign memory[11] = {`ADDI, `ZERO, `T0, 16'd1};
assign memory[12] = {`SW, `SP, `T0, 16'd20};
assign memory[13] = {`ADDI, `ZERO, `T0, 16'd6};
assign memory[14] = {`SW, `SP, `T0, 16'd24};
assign memory[15] = {`LUI, `NULL, `T5, 16'd65535};
assign memory[16] = {`ORI, `T5, `T5, 16'd12};
assign memory[17] = {`ADDI, `ZERO, `S0, 16'd10};
assign memory[18] = {`ADDI, `ZERO, `S1, 16'd10};
assign memory[19] = {`ADDI, `ZERO, `S2, 16'd1};
assign memory[20] = {`ADDI, `ZERO, `S3, -16'd1};
assign memory[21] = {`LUI, `NULL, `A0, 16'd4};
assign memory[22] = {`SPECIAL, `ZERO, `S0, `T7, 5'd0, `ADD};
assign memory[23] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[24] = {`SPECIAL, `T7, `S1, `T7, 5'd0, `OR};
assign memory[25] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[26] = {`SW, `T5, `A0, 16'd0};
assign memory[27] = {`ADDI, `ZERO, `S4, 16'd2};
assign memory[28] = {`ADDI, `ZERO, `S5, 16'd5};
assign memory[29] = {`LW, `SP, `T0, 16'd24};
assign memory[30] = {`SPECIAL, `NULL, `T0, `T1, 5'd1, `SRA};
assign memory[31] = {`SPECIAL, `S1, `ZERO, `S5, 5'd0, `ADD};
assign memory[32] = {`LUI, `NULL, `A0, 16'd2};
assign memory[33] = {`SPECIAL, `ZERO, `S4, `T7, 5'd0, `ADD};
assign memory[34] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[35] = {`SPECIAL, `T7, `S5, `T7, 5'd0, `OR};
assign memory[36] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[37] = {`SW, `T5, `A0, 16'd0};
assign memory[38] = {`LUI, `NULL, `A0, 16'd2};
assign memory[39] = {`SPECIAL, `ZERO, `S4, `T7, 5'd0, `ADD};
assign memory[40] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[41] = {`ADDI, `T1, `T2, -16'd1};
assign memory[42] = {`SPECIAL, `S5, `T2, `T6, 5'd0, `SUB};
assign memory[43] = {`SPECIAL, `T7, `T6, `T7, 5'd0, `OR};
assign memory[44] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[45] = {`SW, `T5, `A0, 16'd0};
assign memory[46] = {`ADDI, `T1, `T1, -16'd1};
assign memory[47] = {`BNE, `T1, `ZERO, -16'd16};
assign memory[48] = {`NOP};
assign memory[49] = {`ADDI, `SP, `SP, -16'd4};
assign memory[50] = {`SW, `SP, `RA, 16'd0};
assign memory[51] = {`JAL, 26'd86};
assign memory[52] = {`NOP};
assign memory[53] = {`LW, `SP, `RA, 16'd0};
assign memory[54] = {`ADDI, `SP, `SP, 16'd4};
assign memory[55] = {`ADDI, `ZERO, `T0, 16'd1};
assign memory[56] = {`SPECIAL, `T0, `S1, `T0, 5'd0, `SLT};
assign memory[57] = {`BEQ, `T0, `ZERO, 16'd8};
assign memory[58] = {`NOP};
assign memory[59] = {`ADDI, `ZERO, `T0, 16'd27};
assign memory[60] = {`SPECIAL, `S1, `T0, `T0, 5'd0, `SLT};
assign memory[61] = {`BEQ, `T0, `ZERO, 16'd5};
assign memory[62] = {`NOP};
assign memory[63] = {`ADDI, `SP, `SP, -16'd4};
assign memory[64] = {`SW, `SP, `RA, 16'd0};
assign memory[65] = {`JAL, 26'd105};
assign memory[66] = {`NOP};
assign memory[67] = {`LW, `SP, `RA, 16'd0};
assign memory[68] = {`ADDI, `SP, `SP, 16'd4};
assign memory[69] = {`ADDI, `ZERO, `T1, 16'd32767};
assign memory[70] = {`ADDI, `T1, `T1, -16'd1};
assign memory[71] = {`BNE, `T1, `ZERO, -16'd2};
assign memory[72] = {`NOP};
assign memory[73] = {`SPECIAL, `ZERO, `ZERO, `T1, 5'd0, `ADD};
assign memory[74] = {`LW, `SP, `T0, 16'd0};
assign memory[75] = {`SPECIAL, `S0, `T0, `T4, 5'd0, `SLT};
assign memory[76] = {`BEQ, `T4, `ZERO, 16'd74};
assign memory[77] = {`NOP};
assign memory[78] = {`LW, `SP, `T0, 16'd4};
assign memory[79] = {`SPECIAL, `S1, `T0, `T4, 5'd0, `SLT};
assign memory[80] = {`BEQ, `T4, `ZERO, 16'd75};
assign memory[81] = {`NOP};
assign memory[82] = {`ADDI, `T1, `T1, 16'd1};
assign memory[83] = {`SPECIAL, `ZERO, `ZERO, `T0, 5'd0, `ADD};
assign memory[84] = {`SPECIAL, `T0, `S1, `T4, 5'd0, `SLT};
assign memory[85] = {`BEQ, `T4, `ZERO, 16'd71};
assign memory[86] = {`NOP};
assign memory[87] = {`SPECIAL, `T0, `S0, `T4, 5'd0, `SLT};
assign memory[88] = {`BEQ, `T4, `ZERO, 16'd3};
assign memory[89] = {`NOP};
assign memory[90] = {`ADDI, `S4, `T0, 16'd1};
assign memory[91] = {`BEQ, `S0, `T0, 16'd71};
assign memory[92] = {`NOP};
assign memory[93] = {`J, 26'd48};
assign memory[94] = {`NOP};
assign memory[95] = {`ADDI, `ZERO, `A0, 16'd69};
assign memory[96] = {`SW, `T5, `A0, 16'd0};
assign memory[97] = {`ADDI, `ZERO, `V0, 16'd10};
assign memory[98] = {`ADDI, `SP, `SP, -16'd4};
assign memory[99] = {`SW, `SP, `RA, 16'd0};
assign memory[100] = {`LUI, `NULL, `A0, 16'd0};
assign memory[101] = {`SPECIAL, `ZERO, `S0, `T7, 5'd0, `ADD};
assign memory[102] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[103] = {`SPECIAL, `T7, `S1, `T7, 5'd0, `OR};
assign memory[104] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[105] = {`SW, `T5, `A0, 16'd0};
assign memory[106] = {`SPECIAL, `S0, `S2, `S0, 5'd0, `ADD};
assign memory[107] = {`SPECIAL, `S1, `S3, `S1, 5'd0, `ADD};
assign memory[108] = {`LUI, `NULL, `A0, 16'd4};
assign memory[109] = {`SPECIAL, `ZERO, `S0, `T7, 5'd0, `ADD};
assign memory[110] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[111] = {`SPECIAL, `T7, `S1, `T7, 5'd0, `OR};
assign memory[112] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[113] = {`SW, `T5, `A0, 16'd0};
assign memory[114] = {`LW, `SP, `RA, 16'd0};
assign memory[115] = {`ADDI, `SP, `SP, 16'd4};
assign memory[116] = {`SPECIAL, `RA, `NULL, `NULL, 5'd0, `JR};
assign memory[117] = {`NOP};
assign memory[118] = {`LW, `SP, `T0, 16'd28};
assign memory[119] = {`SPECIAL, `NULL, `T0, `T1, 5'd1, `SRA};
assign memory[120] = {`ADDI, `SP, `SP, -16'd4};
assign memory[121] = {`SW, `SP, `RA, 16'd0};
assign memory[122] = {`SPECIAL, `S3, `ZERO, `T2, 5'd0, `SLT};
assign memory[123] = {`BEQ, `T2, `ZERO, 16'd16};
assign memory[124] = {`NOP};
assign memory[125] = {`ADDI, `S5, `T2, 16'd3};
assign memory[126] = {`LUI, `NULL, `A0, 16'd0};
assign memory[127] = {`SPECIAL, `ZERO, `S4, `T7, 5'd0, `ADD};
assign memory[128] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[129] = {`SPECIAL, `T7, `T2, `T7, 5'd0, `OR};
assign memory[130] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[131] = {`SW, `T5, `A0, 16'd0};
assign memory[132] = {`ADDI, `S5, `T2, -16'd3};
assign memory[133] = {`LUI, `NULL, `A0, 16'd2};
assign memory[134] = {`SPECIAL, `ZERO, `S4, `T7, 5'd0, `ADD};
assign memory[135] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[136] = {`SPECIAL, `T7, `T2, `T7, 5'd0, `OR};
assign memory[137] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[138] = {`SW, `T5, `A0, 16'd0};
assign memory[139] = {`SPECIAL, `S1, `ZERO, `S5, 5'd0, `ADD};
assign memory[140] = {`J, 26'd142};
assign memory[141] = {`NOP};
assign memory[142] = {`ADDI, `S5, `T2, -16'd2};
assign memory[143] = {`LUI, `NULL, `A0, 16'd0};
assign memory[144] = {`SPECIAL, `ZERO, `S4, `T7, 5'd0, `ADD};
assign memory[145] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[146] = {`SPECIAL, `T7, `T2, `T7, 5'd0, `OR};
assign memory[147] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[148] = {`SW, `T5, `A0, 16'd0};
assign memory[149] = {`ADDI, `S5, `T2, 16'd4};
assign memory[150] = {`LUI, `NULL, `A0, 16'd2};
assign memory[151] = {`SPECIAL, `ZERO, `S4, `T7, 5'd0, `ADD};
assign memory[152] = {`SPECIAL, `NULL, `T7, `T7, 5'd8, `SLL};
assign memory[153] = {`SPECIAL, `T7, `T2, `T7, 5'd0, `OR};
assign memory[154] = {`SPECIAL, `A0, `T7, `A0, 5'd0, `OR};
assign memory[155] = {`SW, `T5, `A0, 16'd0};
assign memory[156] = {`SPECIAL, `S1, `ZERO, `S5, 5'd0, `ADD};
assign memory[157] = {`LW, `SP, `RA, 16'd0};
assign memory[158] = {`ADDI, `SP, `SP, 16'd4};
assign memory[159] = {`SPECIAL, `RA, `NULL, `NULL, 5'd0, `JR};
assign memory[160] = {`NOP};
assign memory[161] = {`SPECIAL, `S2, `ZERO, `S2, 5'd0, `NOR};
assign memory[162] = {`ADDI, `S2, `S2, 16'd1};
assign memory[163] = {`BEQ, `T1, `ZERO, -16'd77};
assign memory[164] = {`NOP};
assign memory[165] = {`J, 26'd82};
assign memory[166] = {`NOP};
assign memory[167] = {`SPECIAL, `S3, `ZERO, `S3, 5'd0, `NOR};
assign memory[168] = {`ADDI, `S3, `S3, 16'd1};
assign memory[169] = {`BEQ, `T1, `ZERO, -16'd78};
assign memory[170] = {`NOP};
assign memory[171] = {`J, 26'd78};
assign memory[172] = {`NOP};
assign memory[173] = {`ADDI, `S5, `T2, -16'd2};
assign memory[174] = {`SPECIAL, `T2, `S1, `T3, 5'd0, `SLT};
assign memory[175] = {`BEQ, `T3, `ZERO, 16'd4};
assign memory[176] = {`NOP};
assign memory[177] = {`ADDI, `S5, `T2, 16'd3};
assign memory[178] = {`SPECIAL, `S1, `T2, `T3, 5'd0, `SLT};
assign memory[179] = {`BEQ, `T3, `ZERO, 16'd1};
assign memory[180] = {`NOP};
assign memory[181] = {`J, 26'd145};
assign memory[182] = {`NOP};
assign memory[183] = {`J, 26'd82};
    assign memory[184] = {`NOP};
    assign memory[185] = {`NOP};
    assign memory[186] = {`NOP};
    assign memory[187] = {`NOP};
    assign memory[188] = {`NOP};
    assign memory[189] = {`NOP};
    assign memory[190] = {`NOP};
    assign memory[191] = {`NOP};
    assign memory[192] = {`NOP};
    assign memory[193] = {`NOP};
    assign memory[194] = {`NOP};
    assign memory[195] = {`NOP};
    assign memory[196] = {`NOP};
    assign memory[197] = {`NOP};
    assign memory[198] = {`NOP};
    assign memory[199] = {`NOP};
    assign memory[200] = {`NOP};
    assign memory[201] = {`NOP};
    assign memory[202] = {`NOP};
    assign memory[203] = {`NOP};
    assign memory[204] = {`NOP};
    assign memory[205] = {`NOP};
    assign memory[206] = {`NOP};
    assign memory[207] = {`NOP};
    assign memory[208] = {`NOP};
    assign memory[209] = {`NOP};
    assign memory[210] = {`NOP};
    assign memory[211] = {`NOP};
    assign memory[212] = {`NOP};
    assign memory[213] = {`NOP};
    assign memory[214] = {`NOP};
    assign memory[215] = {`NOP};
    assign memory[216] = {`NOP};
    assign memory[217] = {`NOP};
    assign memory[218] = {`NOP};
    assign memory[219] = {`NOP};
    assign memory[220] = {`NOP};
    assign memory[221] = {`NOP};
    assign memory[222] = {`NOP};
    assign memory[223] = {`NOP};
    assign memory[224] = {`NOP};
    assign memory[225] = {`NOP};
    assign memory[226] = {`NOP};
    assign memory[227] = {`NOP};
    assign memory[228] = {`NOP};
    assign memory[229] = {`NOP};
    assign memory[230] = {`NOP};
    assign memory[231] = {`NOP};
    assign memory[232] = {`NOP};
    assign memory[233] = {`NOP};
    assign memory[234] = {`NOP};
    assign memory[235] = {`NOP};
    assign memory[236] = {`NOP};
    assign memory[237] = {`NOP};
    assign memory[238] = {`NOP};
    assign memory[239] = {`NOP};
    assign memory[240] = {`NOP};
    assign memory[241] = {`NOP};
    assign memory[242] = {`NOP};
    assign memory[243] = {`NOP};
    assign memory[244] = {`NOP};
    assign memory[245] = {`NOP};
    assign memory[246] = {`NOP};
    assign memory[247] = {`NOP};
    assign memory[248] = {`NOP};
    assign memory[249] = {`NOP};
    assign memory[250] = {`NOP};
    assign memory[251] = {`NOP};
    assign memory[252] = {`NOP};
    assign memory[253] = {`NOP};
    assign memory[254] = {`NOP};
    assign memory[255] = {`NOP};
    assign memory[256] = {`NOP};
    assign memory[257] = {`NOP};
    assign memory[258] = {`NOP};
    assign memory[259] = {`NOP};
    assign memory[260] = {`NOP};
    assign memory[261] = {`NOP};
    assign memory[262] = {`NOP};
    assign memory[263] = {`NOP};
    assign memory[264] = {`NOP};
    assign memory[265] = {`NOP};
    assign memory[266] = {`NOP};
    assign memory[267] = {`NOP};
    assign memory[268] = {`NOP};
    assign memory[269] = {`NOP};
    assign memory[270] = {`NOP};
    assign memory[271] = {`NOP};
    assign memory[272] = {`NOP};
    assign memory[273] = {`NOP};
    assign memory[274] = {`NOP};
    assign memory[275] = {`NOP};
    assign memory[276] = {`NOP};
    assign memory[277] = {`NOP};
    assign memory[278] = {`NOP};
    assign memory[279] = {`NOP};
    assign memory[280] = {`NOP};
    assign memory[281] = {`NOP};
    assign memory[282] = {`NOP};
    assign memory[283] = {`NOP};
    assign memory[284] = {`NOP};
    assign memory[285] = {`NOP};
    assign memory[286] = {`NOP};
    assign memory[287] = {`NOP};
    assign memory[288] = {`NOP};
    assign memory[289] = {`NOP};
    assign memory[290] = {`NOP};
    assign memory[291] = {`NOP};
    assign memory[292] = {`NOP};
    assign memory[293] = {`NOP};
    assign memory[294] = {`NOP};
    assign memory[295] = {`NOP};
    assign memory[296] = {`NOP};
    assign memory[297] = {`NOP};
    assign memory[298] = {`NOP};
    assign memory[299] = {`NOP};
    assign memory[300] = {`NOP};
    assign memory[301] = {`NOP};
    assign memory[302] = {`NOP};
    assign memory[303] = {`NOP};
    assign memory[304] = {`NOP};
    assign memory[305] = {`NOP};
    assign memory[306] = {`NOP};
    assign memory[307] = {`NOP};
    assign memory[308] = {`NOP};
    assign memory[309] = {`NOP};
    assign memory[310] = {`NOP};
    assign memory[311] = {`NOP};
    assign memory[312] = {`NOP};
    assign memory[313] = {`NOP};
    assign memory[314] = {`NOP};
    assign memory[315] = {`NOP};
    assign memory[316] = {`NOP};
    assign memory[317] = {`NOP};
    assign memory[318] = {`NOP};
    assign memory[319] = {`NOP};
    assign memory[320] = {`NOP};
    assign memory[321] = {`NOP};
    assign memory[322] = {`NOP};
    assign memory[323] = {`NOP};
    assign memory[324] = {`NOP};
    assign memory[325] = {`NOP};
    assign memory[326] = {`NOP};
    assign memory[327] = {`NOP};
    assign memory[328] = {`NOP};
    assign memory[329] = {`NOP};
    assign memory[330] = {`NOP};
    assign memory[331] = {`NOP};
    assign memory[332] = {`NOP};
    assign memory[333] = {`NOP};
    assign memory[334] = {`NOP};
    assign memory[335] = {`NOP};
    assign memory[336] = {`NOP};
    assign memory[337] = {`NOP};
    assign memory[338] = {`NOP};
    assign memory[339] = {`NOP};
    assign memory[340] = {`NOP};
    assign memory[341] = {`NOP};
    assign memory[342] = {`NOP};
    assign memory[343] = {`NOP};
    assign memory[344] = {`NOP};
    assign memory[345] = {`NOP};
    assign memory[346] = {`NOP};
    assign memory[347] = {`NOP};
    assign memory[348] = {`NOP};
    assign memory[349] = {`NOP};
    assign memory[350] = {`NOP};
    assign memory[351] = {`NOP};
    assign memory[352] = {`NOP};
    assign memory[353] = {`NOP};
    assign memory[354] = {`NOP};
    assign memory[355] = {`NOP};
    assign memory[356] = {`NOP};
    assign memory[357] = {`NOP};
    assign memory[358] = {`NOP};
    assign memory[359] = {`NOP};
    assign memory[360] = {`NOP};
    assign memory[361] = {`NOP};
    assign memory[362] = {`NOP};
    assign memory[363] = {`NOP};
    assign memory[364] = {`NOP};
    assign memory[365] = {`NOP};
    assign memory[366] = {`NOP};
    assign memory[367] = {`NOP};
    assign memory[368] = {`NOP};
    assign memory[369] = {`NOP};
    assign memory[370] = {`NOP};
    assign memory[371] = {`NOP};
    assign memory[372] = {`NOP};
    assign memory[373] = {`NOP};
    assign memory[374] = {`NOP};
    assign memory[375] = {`NOP};
    assign memory[376] = {`NOP};
    assign memory[377] = {`NOP};
    assign memory[378] = {`NOP};
    assign memory[379] = {`NOP};
    assign memory[380] = {`NOP};
    assign memory[381] = {`NOP};
    assign memory[382] = {`NOP};
    assign memory[383] = {`NOP};
    assign memory[384] = {`NOP};
    assign memory[385] = {`NOP};
    assign memory[386] = {`NOP};
    assign memory[387] = {`NOP};
    assign memory[388] = {`NOP};
    assign memory[389] = {`NOP};
    assign memory[390] = {`NOP};
    assign memory[391] = {`NOP};
    assign memory[392] = {`NOP};
    assign memory[393] = {`NOP};
    assign memory[394] = {`NOP};
    assign memory[395] = {`NOP};
    assign memory[396] = {`NOP};
    assign memory[397] = {`NOP};
    assign memory[398] = {`NOP};
    assign memory[399] = {`NOP};
    assign memory[400] = {`NOP};
    assign memory[401] = {`NOP};
    assign memory[402] = {`NOP};
    assign memory[403] = {`NOP};
    assign memory[404] = {`NOP};
    assign memory[405] = {`NOP};
    assign memory[406] = {`NOP};
    assign memory[407] = {`NOP};
    assign memory[408] = {`NOP};
    assign memory[409] = {`NOP};
    assign memory[410] = {`NOP};
    assign memory[411] = {`NOP};
    assign memory[412] = {`NOP};
    assign memory[413] = {`NOP};
    assign memory[414] = {`NOP};
    assign memory[415] = {`NOP};
    assign memory[416] = {`NOP};
    assign memory[417] = {`NOP};
    assign memory[418] = {`NOP};
    assign memory[419] = {`NOP};
    assign memory[420] = {`NOP};
    assign memory[421] = {`NOP};
    assign memory[422] = {`NOP};
    assign memory[423] = {`NOP};
    assign memory[424] = {`NOP};
    assign memory[425] = {`NOP};
    assign memory[426] = {`NOP};
    assign memory[427] = {`NOP};
    assign memory[428] = {`NOP};
    assign memory[429] = {`NOP};
    assign memory[430] = {`NOP};
    assign memory[431] = {`NOP};
    assign memory[432] = {`NOP};
    assign memory[433] = {`NOP};
    assign memory[434] = {`NOP};
    assign memory[435] = {`NOP};
    assign memory[436] = {`NOP};
    assign memory[437] = {`NOP};
    assign memory[438] = {`NOP};
    assign memory[439] = {`NOP};
    assign memory[440] = {`NOP};
    assign memory[441] = {`NOP};
    assign memory[442] = {`NOP};
    assign memory[443] = {`NOP};
    assign memory[444] = {`NOP};
    assign memory[445] = {`NOP};
    assign memory[446] = {`NOP};
    assign memory[447] = {`NOP};
    assign memory[448] = {`NOP};
    assign memory[449] = {`NOP};
    assign memory[450] = {`NOP};
    assign memory[451] = {`NOP};
    assign memory[452] = {`NOP};
    assign memory[453] = {`NOP};
    assign memory[454] = {`NOP};
    assign memory[455] = {`NOP};
    assign memory[456] = {`NOP};
    assign memory[457] = {`NOP};
    assign memory[458] = {`NOP};
    assign memory[459] = {`NOP};
    assign memory[460] = {`NOP};
    assign memory[461] = {`NOP};
    assign memory[462] = {`NOP};
    assign memory[463] = {`NOP};
    assign memory[464] = {`NOP};
    assign memory[465] = {`NOP};
    assign memory[466] = {`NOP};
    assign memory[467] = {`NOP};
    assign memory[468] = {`NOP};
    assign memory[469] = {`NOP};
    assign memory[470] = {`NOP};
    assign memory[471] = {`NOP};
    assign memory[472] = {`NOP};
    assign memory[473] = {`NOP};
    assign memory[474] = {`NOP};
    assign memory[475] = {`NOP};
    assign memory[476] = {`NOP};
    assign memory[477] = {`NOP};
    assign memory[478] = {`NOP};
    assign memory[479] = {`NOP};
    assign memory[480] = {`NOP};
    assign memory[481] = {`NOP};
    assign memory[482] = {`NOP};
    assign memory[483] = {`NOP};
    assign memory[484] = {`NOP};
    assign memory[485] = {`NOP};
    assign memory[486] = {`NOP};
    assign memory[487] = {`NOP};
    assign memory[488] = {`NOP};
    assign memory[489] = {`NOP};
    assign memory[490] = {`NOP};
    assign memory[491] = {`NOP};
    assign memory[492] = {`NOP};
    assign memory[493] = {`NOP};
    assign memory[494] = {`NOP};
    assign memory[495] = {`NOP};
    assign memory[496] = {`NOP};
    assign memory[497] = {`NOP};
    assign memory[498] = {`NOP};
    assign memory[499] = {`NOP};
    assign memory[500] = {`NOP};
    assign memory[501] = {`NOP};
    assign memory[502] = {`NOP};
    assign memory[503] = {`NOP};
    assign memory[504] = {`NOP};
    assign memory[505] = {`NOP};
    assign memory[506] = {`NOP};
    assign memory[507] = {`NOP};
    assign memory[508] = {`NOP};
    assign memory[509] = {`NOP};
    assign memory[510] = {`NOP};
    assign memory[511] = {`NOP};

endmodule
