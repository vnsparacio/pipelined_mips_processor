`include "mips_defines.v"

`define ADDR_WIDTH 9
`define INSTR_WIDTH 32
`define NUM_INSTR 512

module pong_irom_VS(clk, addr, dout);
    input clk;
    input [`ADDR_WIDTH-1:0] addr;
    output reg [`INSTR_WIDTH-1:0] dout;
    
    wire [`INSTR_WIDTH-1:0] memory [`NUM_INSTR-1:0];
    
    always @(posedge clk)
        dout <= memory[addr];

    // without forwarding, we need two cycles of NOPs before
    // data can be used
    // implement lots of tests here, and make another irom.v
    // with your implementation of Pong
    // don't forget that this processor has a branch delay slot
    assign memory[  0] = {`LUI, `NULL, `T0, 16'hffff};
    assign memory[  1] = {`NOP};
    assign memory[  2] = {`NOP};
    assign memory[  3] = {`ORI, `T0, `T0, 16'h000c};
    assign memory[  4] = {`LUI, `NULL, `T1, 16'h6};
    assign memory[  5] = {`NOP};
    assign memory[  6] = {`ORI, `T1, `T1, 8'd1, 8'd1};
    assign memory[  7] = {`SW, `T0, `T1, 16'd0}; // draws yellow at (1,1)
  assign memory[  8] = {`NOP};
  assign memory[  9] = {`NOP};
  assign memory[ 10] = {`NOP};
  assign memory[ 11] = {`ADDI, `ZERO, `SP, 16'd0}; 
  assign memory[ 12] = {`ADDI, `ZERO, `T0, 16'd39}; //maximum x coordinate
  assign memory[ 13] = {`SW,`SP, `T0,  16'd0};
  assign memory[ 14] = {`ADDI, `ZERO, `T0, 16'd29}; //maximum y  coordinate 
  assign memory[ 15] = {`SW, `SP,`T0,  16'd4};
  assign memory[ 16] = {`ADDI, `ZERO, `T0, 16'd0}; // background color
  assign memory[ 17] = {`SW, `SP,`T0,  16'd8};
  assign memory[ 18] = {`ADDI, `ZERO, `T0, 16'd2}; // paddle color
  assign memory[ 19] = {`SW,`SP, `T0,  16'd12};
  assign memory[ 20] = {`ADDI, `ZERO, `T0, 16'd4}; // ball color
  assign memory[ 21] = {`SW, `SP, `T0,  16'd16};
  assign memory[ 22] = {`ADDI, `ZERO, `T0, 16'd1}; // ball height and width and paddle width 
  assign memory[ 23] = {`SW,`SP,  `T0, 16'd20};
  assign memory[ 24] = {`ADDI, `ZERO, `T0, 16'd6}; // paddle height
  assign memory[ 25] = {`SW,`SP, `T0,  16'd24};
  assign memory[ 26] = {`ADDI, `ZERO, `T0, 16'd1}; // init x coord
  assign memory[ 27] = {`SW, `SP, `T0,  16'd28};    
  assign memory[ 28] = {`ADDI, `ZERO, `T0, 16'd15}; // init y coord
  assign memory[ 29] = {`SW,`SP, `T0,  16'd32}; 
  assign memory[ 30] = {`NOP};
  assign memory[ 31] = {`NOP};
  assign memory[ 32] = {`NOP};
  assign memory[ 33] = {`NOP};
  assign memory[ 34] = {`NOP};
  assign memory[ 35] = {`ADDI, `ZERO, `A0, 16'd0}; // init
  assign memory[ 36] = {`ADDI, `ZERO, `A1, 16'd12};
  assign memory[ 37] = {`ADDI, `ZERO, `A2, 16'd2};
  assign memory[ 38] = {`JAL, 26'd343}; //jump to draw_block
  assign memory[ 39] = {`NOP};
  assign memory[ 40] = {`ADDI, `ZERO, `A0, 16'd39}; 
  assign memory[ 41] = {`ADDI, `ZERO, `A1, 16'd12}; 
  assign memory[ 42] = {`ADDI, `ZERO, `A2, 16'd2}; 
  assign memory[ 43] = {`JAL, 26'd343}; //jump to draw_block
  assign memory[ 44] = {`NOP};
  assign memory[ 45] = {`ADDI, `ZERO, `T4, 16'd1}; //x coordinate  
  assign memory[ 46] = {`NOP}; //{`JAL, 26'd418}; //jump to write_byte
  assign memory[ 47] = {`NOP};
  assign memory[ 48] = {`ADDI, `ZERO, `T5, 16'd15};  //y coordinate
  assign memory[ 49] = {`ADDI, `ZERO, `A0, 16'd1}; //color //{`JAL, 26'd418}; //jump to write_byte
  assign memory[ 50] = {`SPECIAL, `NULL, `A0, `A0, 5'd16, `SLL};
  assign memory[ 51] = {`ORI, `A0, `A0, `T4, `T5}; 
  assign memory[ 52] = {`JAL, 26'd418}; //jump to write_byte
  assign memory[ 53] = {`NOP};
  assign memory[ 54] = {`JAL, 26'd390}; //jump to pause
  assign memory[ 55] = {`NOP}; 
  assign memory[ 56] = {`ADDI, `ZERO, `A0, 16'd0};  
  assign memory[ 57] = {`ADDI, `ZERO, `A1, 16'd12};  
  assign memory[ 58] = {`ADDI, `ZERO, `A2, -16'd1};  
  assign memory[ 59] = {`JAL, 26'd270}; //jump to move_paddle
  assign memory[ 60] = {`NOP}; 

  // game_loop
  assign memory[ 61] = {`ADDI, `ZERO, `T0, 16'd1}; //dX 
  assign memory[ 62] = {`SW, `SP, `T0, 16'd36};
  assign memory[ 63] = {`ADDI, `ZERO, `T0, 16'd1}; //dY: should be able to comment this line out?
  assign memory[ 64] = {`SW, `SP,`T0,  16'd40};
  assign memory[ 65] = {`ADDI, `ZERO, `T0, 16'd12}; //Y coordinate of top of paddle
  assign memory[ 66] = {`SW,`SP, `T0,  16'd44};
  assign memory[ 67] = {`JAL, 26'd138}; //jump to ball_loop_condition
  assign memory[ 68] = {`NOP};
  assign memory[ 69] = {`NOP};
  assign memory[ 70] = {`NOP};
  assign memory[ 71] = {`NOP}; // ball_loop_body
  assign memory[ 72] = {`LW, `SP,`A0,  16'd28};
  assign memory[ 73] = {`LW,`SP, `A1,  16'd32};
  assign memory[ 74] = {`LW, `SP, `A2, 16'd36};
  assign memory[ 75] = {`LW, `SP, `A3, 16'd40};
  assign memory[ 76] = {`JAL, 26'd238}; // jump to move_ball
  assign memory[ 77] = {`NOP};
  assign memory[ 78] = {`JAL, 26'd390}; // jump to pause
  assign memory[ 79] = {`NOP};
  assign memory[ 80] = {`SW,`SP, `V0,  16'd28};
  assign memory[ 81] = {`SW, `SP,`V1,  16'd32};
  assign memory[ 82] = {`LW, `SP,`T0,  16'd44};
  assign memory[ 83] = {`ADDI, `T0, `T0, 16'd3}; 
  assign memory[ 84] = {`SPECIAL, `T0, `V1, `T3, `NULL, `SUB};
  assign memory[ 85] = {`SPECIAL, `T3, `ZERO, `T4, `NULL, `SLT};
  assign memory[ 86] = {`BNE, `T4, `ZERO, 16'ha}; // branch to paddle_move_down
  assign memory[ 87] = {`J, 26'd106};  //jump to paddle_move_up
  assign memory[ 88] = {`NOP};
  assign memory[ 89] = {`NOP};
  assign memory[ 90] = {`NOP}; // paddle_move_down
  assign memory[ 91] = {`ADDI, `T0, `ZERO, 16'd24}; 
  assign memory[ 92] = {`LW, `SP,`A1,  16'd44}; //a1 = t0 = ycoord of top of paddle + 3 = ycoord of "center" of paddle
  assign memory[ 93] = {`SPECIAL, `A1, `T0, `T1, `NULL, `SLT};
  assign memory[ 94] = {`BEQ, `T1, `ZERO, 16'd333}; // paddle_move_skip 
  assign memory[ 95] = {`ADDI, `ZERO, `A2, 16'd0};  // load 0 into A0
  assign memory[ 96] = {`JAL, 26'd270}; // jump to move_paddle
  assign memory[ 97] = {`NOP};
  assign memory[ 98] = {`ADDI, `ZERO, `A0, 16'd39};  
  assign memory[ 99] = {`JAL, 26'd270}; // jump to move_paddle
  assign memory[100] = {`NOP};
  assign memory[101] = {`JAL, 26'd390}; // jump to pause
  assign memory[102] = {`NOP};
  assign memory[103] = {`SW,`SP, `V0,  16'd44};
  assign memory[104] = {`J, 26'd138};  //jump to ball_loop_condition
  assign memory[105] = {`NOP};
  assign memory[106] = {`NOP}; // paddle_move_up
  assign memory[107] = {`ADDI, `ZERO, `T0, 16'd0};  
  assign memory[108] = {`LW, `SP,`A1,  16'd44}; // a1 = t0 = ycoord of top of paddle + 3 = ycoord of "center" of paddle
  assign memory[109] = {`SPECIAL, `T0, `A1, `T1, `NULL, `SLT}; // 0 < A1
  assign memory[110] = {`BEQ, `T1, `ZERO, 16'd19}; // paddle_move_skip 
  assign memory[111] = {`NOP};
  assign memory[112] = {`ADDI, `ZERO, `A0, 16'd0};  
  assign memory[113] = {`ADDI, `ZERO, `A2, -16'd1};  
  assign memory[114] = {`JAL, 26'd270}; // jump to move_paddle
  assign memory[115] = {`NOP};
  assign memory[116] = {`ADDI, `ZERO, `A0, 16'd39};  
  assign memory[117] = {`JAL, 26'd270}; // jump to move_paddle
  assign memory[118] = {`NOP};
  assign memory[119] = {`JAL, 26'd390}; // jump to pause
  assign memory[120] = {`NOP};
  assign memory[121] = {`SW, `SP,`V0,  16'd44};
  assign memory[122] = {`J, 26'd138};  //jump to ball_loop_condition
  assign memory[123] = {`NOP};
  assign memory[124] = {`NOP};
  assign memory[125] = {`NOP};
  assign memory[126] = {`NOP};
  assign memory[127] = {`NOP};
  assign memory[128] = {`NOP};
  assign memory[129] = {`NOP}; // paddle_move_skip
  assign memory[130] = {`JAL, 26'd390}; // jump to pause
  assign memory[131] = {`NOP};
  assign memory[132] = {`J, 26'd138};  //jump to ball_loop_condition
  assign memory[133] = {`NOP};
  assign memory[134] = {`NOP};
  assign memory[135] = {`NOP};
  assign memory[136] = {`NOP};
  assign memory[137] = {`NOP};
  assign memory[138] = {`NOP}; // ball_loop_condition
  assign memory[139] = {`LW, `SP, `T6,  16'd28};
  assign memory[140] = {`ADDI, `ZERO, `T7, 16'd0};
  assign memory[141] = {`BEQ, `T6, `T7, 16'd298}; //end the game 
  assign memory[142] = {`NOP};
  assign memory[143] = {`LW,`SP,  `T6, 16'd28};
  assign memory[144] = {`ADDI, `ZERO, `T7, 16'd39};
  assign memory[145] = {`BEQ, `T6, `T7, 16'd293}; //end the game 
  assign memory[146] = {`NOP};
  assign memory[147] = {`LW, `SP,`T6,  16'd28};
  assign memory[148] = {`ADDI, `ZERO, `T7, 16'd1};
  assign memory[149] = {`SPECIAL, `T6, `T7, `T5, `NULL, `SUB}; //t5 = 0 if xcoord of ball = 1
  assign memory[150] = {`BNE, `T5, `ZERO, 16'ha}; //other_paddle
  assign memory[151] = {`NOP};
  assign memory[152] = {`LW, `SP,`T4,  16'd32}; //ycoordinate of the ball
  assign memory[153] = {`LW, `SP,`T3,  16'd44}; //ycoordinate of the the top of the paddle = t3
  assign memory[154] = {`SPECIAL, `T4, `T3, `T2, `NULL, `SUB}; // t2 = ycoord of ball - ycoord of top of paddle: if t2<0, not within paddle length
  assign memory[155] = {`SPECIAL, `T2, `ZERO, `T1, `NULL, `SLT};
  assign memory[156] = {`BNE, `T1, `ZERO, 16'ha}; //other_paddle
  assign memory[157] = {`NOP};
  assign memory[158] = {`ADDI, `ZERO, `T1, 16'd6};
  assign memory[159] = {`SPECIAL, `T2, `T1, `T0, `NULL, `SLT}; //ycoord of bal-ycoord of paddle< 6
  assign memory[160] = {`BEQ, `T0, `ZERO, 16'd9}; //other_paddle 
  assign memory[161] = {`NOP};
  assign memory[162] = {`ADDI, `ZERO, `T0, 16'd1};
  assign memory[163] = {`SW, `SP, `T0,  16'd36};
  assign memory[164] = {`NOP};
  assign memory[165] = {`NOP};
  assign memory[166] = {`NOP};
  assign memory[167] = {`NOP};
  assign memory[168] = {`NOP};
  assign memory[169] = {`NOP};//other_paddle
  assign memory[170] = {`LW,`SP, `T6,  16'd28};
  assign memory[171] = {`ADDI, `ZERO, `T7, 16'd38};
  assign memory[172] = {`SPECIAL, `T6, `T7, `T5, `NULL, `SUB}; // #t5 = 0 if xcoord of ball = 38
  assign memory[173] = {`BNE, `T5, `ZERO, 16'd19}; //continue
  assign memory[174] = {`NOP};
  assign memory[175] = {`LW, `SP, `T4,  16'd32}; //ycoord of the ball
  assign memory[176] = {`LW, `SP, `T3,  16'd44}; //t3 = ycoord of top of paddle
  assign memory[177] = {`SPECIAL, `T4, `T3, `T2, `NULL, `SUB}; // t2 = ycoord of ball - ycoord of top of paddle: if t2<0, not within paddle length
  assign memory[178] = {`SPECIAL, `T2, `ZERO, `T1, `NULL, `SLT}; 
  assign memory[179] = {`BNE, `T1, `ZERO, 16'd12}; //if t2<0, continue
  assign memory[180] = {`NOP};
  assign memory[181] = {`ADDI, `ZERO, `T1, 16'd6};
  assign memory[182] = {`SPECIAL, `T2, `T1, `T0, `NULL, `SLT}; // ycoord of bal - ycoord of paddle < 6
  assign memory[183] = {`BEQ, `T0, `ZERO, 16'd8}; //continue 
  assign memory[184] = {`NOP};
  assign memory[185] = {`ADDI, `ZERO, `T0, -16'd1};
  assign memory[186] = {`SW, `SP,`T0,  16'd36};
  assign memory[187] = {`NOP};
  assign memory[188] = {`NOP};
  assign memory[189] = {`NOP};
  assign memory[190] = {`NOP};
  assign memory[191] = {`NOP};
  assign memory[192] = {`NOP}; //continue
  assign memory[193] = {`LW,`SP, `T6,  16'd32};
  assign memory[194] = {`ADDI, `ZERO, `T7, 16'd0};
  assign memory[195] = {`BEQ, `T6, `T7, 16'd23}; //y_top_edge
  assign memory[196] = {`NOP};
  assign memory[197] = {`LW, `SP, `T6,  16'd32}; 
  assign memory[198] = {`ADDI, `ZERO, `T7, 16'd29};
  assign memory[199] = {`BEQ, `T6, `T7, 16'd28}; //y_bottom_edge
  assign memory[200] = {`NOP};
  assign memory[201] = {`J, 26'd71};  //ball_loop_body
  assign memory[202] = {`NOP};
  assign memory[203] = {`NOP};
  assign memory[204] = {`NOP};
  assign memory[205] = {`NOP};
  assign memory[206] = {`NOP};
  assign memory[207] = {`NOP};
  assign memory[208] = {`NOP}; // x_right_edge
  assign memory[209] = {`ADDI, `ZERO, `T0, -16'd1};
  assign memory[210] = {`SW, `SP, `T0,  16'd36};
  assign memory[211] = {`J, 26'd192};  //continue
  assign memory[212] = {`NOP};
  assign memory[213] = {`NOP};
  assign memory[214] = {`NOP};
  assign memory[215] = {`NOP};
  assign memory[216] = {`NOP};
  assign memory[217] = {`NOP};
  assign memory[218] = {`NOP};
  assign memory[219] = {`NOP}; // y_top_edge
  assign memory[220] = {`ADDI, `ZERO, `T0, 16'd1};
  assign memory[221] = {`SW,`SP,  `T0, 16'd40};
  assign memory[222] = {`J, 26'd71};  //ball_loop_body
  assign memory[223] = {`NOP};
  assign memory[224] = {`NOP};
  assign memory[225] = {`NOP};
  assign memory[226] = {`NOP};
  assign memory[227] = {`NOP};
  assign memory[228] = {`NOP}; // y_bottom_edge
  assign memory[229] = {`ADDI, `ZERO, `T0, -16'd1};
  assign memory[230] = {`SW,`SP,  `T0, 16'd40};
  assign memory[231] = {`J, 26'd71};  //ball_loop_body
  assign memory[232] = {`NOP};
  assign memory[233] = {`NOP};
  assign memory[234] = {`NOP};
  assign memory[235] = {`NOP};
  assign memory[236] = {`NOP};
  assign memory[237] = {`NOP}; // Game Code Goes Here
  assign memory[238] = {`NOP};// move_ball
  assign memory[239] = {`ADDI, `SP, `SP, -16'd8}; //draws over old ball
  assign memory[240] = {`SW,`SP,  `A0, 16'd0}; //xcoord
  assign memory[241] = {`SW,`SP, `RA,  16'd4};
  assign memory[242] = {`NOP}; //{`JAL, //write_byte a0 is already the x coord
  assign memory[243] = {`ADDI, `A0, `T4, 16'd0}; //T0 becomes x coordinate
  assign memory[244] = {`SPECIAL, `ZERO, `A1, `T5, `NULL, `ADD};  //T1 is the y coord
  assign memory[245] = {`NOP}; //{`JAL, 26'd418}; //write_byte 
  assign memory[246] = {`ADDI, `ZERO, `A0, 16'd0}; //black write byte is stored in A0
  assign memory[247] = {`SPECIAL, `NULL, `A0, `A0, 5'd16, `SLL};
  assign memory[248] = {`ORI, `A0, `A0, `T4, `T5};
  assign memory[249] = {`JAL, 26'd418}; //write_byte 
  assign memory[250] = {`NOP}; //draw new ball
  assign memory[251] = {`LW,`SP, `A0,  16'd0}; 
  assign memory[252] = {`SPECIAL, `A2, `A0, `T4, `NULL, `ADD}; //x coordinate
  assign memory[253] = {`SPECIAL, `ZERO, `A0, `V0, `NULL, `ADD}; //return the new x coord in v0
  assign memory[254] = {`NOP}; //{`JAL, 26'd418}; //write_byte 
  assign memory[255] = {`NOP};
  assign memory[256] = {`SPECIAL, `A3, `A1, `T5, `NULL, `ADD}; //y coordinate
  assign memory[257] = {`SPECIAL, `ZERO, `A0, `V1, `NULL, `ADD};
  assign memory[258] = {`ADDI, `ZERO, `A0, 16'd1}; //color
  assign memory[259] = {`SPECIAL, `NULL, `A0, `A0, 5'd16, `SLL};
  assign memory[260] = {`ORI, `A0, `A0, `T4, `T5};
  assign memory[261] = {`JAL, 26'd418}; //write_byte
  assign memory[262] = {`NOP};
  assign memory[263] = {`LW,`SP, `A0,  16'd0}; 
  assign memory[264] = {`LW,`SP,  `RA, 16'd4}; 
  assign memory[265] = {`ADDI, `SP, `SP, 16'd8};
  assign memory[266] = {`SPECIAL, `RA, 15'd0, `JR};
  assign memory[267] = {`NOP};
  assign memory[268] = {`NOP};
  assign memory[269] = {`NOP};
  assign memory[270] = {`NOP}; // move_paddle
  assign memory[271] = {`ADDI, `SP, `SP, -16'd16};
  assign memory[272] = {`SW,`SP, `A2,  16'd0};
  assign memory[273] = {`SW,`SP, `A1,  16'd4};
  assign memory[274] = {`SW,`SP, `RA,  16'd8};
  assign memory[275] = {`SW, `SP, `A0, 16'd12};
  assign memory[276] = {`ADDI, `ZERO, `A2, 16'd0};
  assign memory[277] = {`JAL, 26'd343}; //draw_block
  assign memory[278] = {`NOP};
  assign memory[279] = {`SPECIAL, `A1, `A2, `V0, `NULL, `ADD};
  assign memory[280] = {`SPECIAL, `A2, `ZERO, `T0, `NULL, `SLT};
  assign memory[281] = {`BNE, `T0, `ZERO, 16'd6}; //move_up if delta is < 0, i.e. delta = -1, the move paddle up
  assign memory[282] = {`NOP};
  assign memory[283] = {`J, 26'd311}; //move_down
  assign memory[284] = {`NOP};
  assign memory[285] = {`NOP};
  assign memory[286] = {`NOP};
  assign memory[287] = {`NOP}; //move_up
  assign memory[288] = {`ADDI, `A1, `S0, 16'd0}; //x coord is 0 so no need to shift
  assign memory[289] = {`SPECIAL, `NULL, `S0, `S0, 5'd16, `SLL};
  assign memory[290] = {`ADDI, `A1, `T0, 16'd5}; //y coord
  assign memory[291] = {`SPECIAL, `ZERO, `T0, `A0, `NULL, `ADD}; 
  assign memory[292] = {`NOP};//{`JAL, 26'd418}; ///////////////////write_byte
  assign memory[293] = {`NOP};
  assign memory[294] = {`ORI, `T0, `A0, `S0, `A0};
  assign memory[295] = {`JAL, 26'd418}; //write_byte //writes the paddle
  assign memory[296] = {`NOP};
  assign memory[297] = {`LW,`SP, `T0,  16'd12}; 	//x coordinate
  assign memory[298] = {`NOP}; 
  assign memory[299] = {`NOP};
  assign memory[300] = {`LW,`SP,  `T1, 16'd4}; 		//y coordinate
  assign memory[301] = {`ADDI, `T1, `T1, -16'd1};
  assign memory[302] = {`ADDI, `ZERO, `A0, 16'd2}; //green color
  assign memory[303] = {`SPECIAL, `NULL, `A0, `A0, 5'd16, `SLL};
  assign memory[304] = {`ORI, `A0, `A0, `T0, `T1}; //A0 = A0 or'ed with {x, y}
  assign memory[305] = {`JAL, 26'd418}; //write_byte
  assign memory[306] = {`NOP};
  assign memory[307] = {`J, 26'd333};  //end_of_move_paddle
  assign memory[308] = {`NOP};
  assign memory[309] = {`NOP};
  assign memory[310] = {`NOP};
  assign memory[311] = {`NOP}; // move_down
  assign memory[312] = {`LW,`SP, `T0,  16'd12}; 		//x coordinate
  assign memory[313] = {`LW,`SP, `T1,  16'd4}; 			//y coordinate
  assign memory[314] = {`ADDI, `ZERO, `A0, 16'd0}; 		//black color
  assign memory[315] = {`SPECIAL, `NULL, `A0, `A0, 5'd16, `SLL};
  assign memory[316] = {`ORI, `A0, `A0, `T0, `T1};
  assign memory[317] = {`JAL, 26'd418}; //write_byte
  assign memory[318] = {`NOP};
  assign memory[319] = {`NOP};
  assign memory[320] = {`NOP};
  assign memory[321] = {`LW,`SP, `T0,  16'd12}; 		//x coordinate
  assign memory[322] = {`LW, `SP, `T1,  16'd4}; 			
  assign memory[323] = {`ADDI, `T1, `T1, 16'd6}; 		//y coordinate
  assign memory[324] = {`ADDI, `ZERO, `A0, 16'd2}; 		//green color
  assign memory[325] = {`SPECIAL, `NULL, `A0, `A0, 5'd16, `SLL};
  assign memory[326] = {`ORI, `A0, `A0, `T0, `T1};
  assign memory[327] = {`JAL, 26'd418}; //write_byte 
  assign memory[328] = {`NOP};
  assign memory[329] = {`NOP};
  assign memory[330] = {`NOP};
  assign memory[331] = {`NOP};
  assign memory[332] = {`NOP};
  assign memory[333] = {`NOP}; // end_of_move_paddle
  assign memory[334] = {`LW, `SP, `A1, 16'd4}; 
  assign memory[335] = {`LW,`SP, `A2,  16'd0}; 
  assign memory[336] = {`LW,`SP, `A0,  16'd12}; 
  assign memory[337] = {`LW,`SP, `RA,  16'd8}; 
  assign memory[338] = {`ADDI, `SP, `SP, 16'd16};
  assign memory[339] = {`SPECIAL, `RA, 15'd0, `JR};
  assign memory[340] = {`NOP};
  assign memory[341] = {`NOP};
  assign memory[342] = {`NOP};//{`SPECIAL, `NULL, `T0, `T0, 5'd16, `SLL}; I have no idea what this is?
  assign memory[343] = {`NOP}; // draw_block
  assign memory[344] = {`ADDI, `SP, `SP, -16'd32};
  assign memory[345] = {`SW,`SP, `A0,  16'd0};
  assign memory[346] = {`SW,`SP, `A1,  16'd4};
  assign memory[347] = {`SW, `SP, `A2, 16'd8};
  assign memory[348] = {`SW, `SP, `A0, 16'd12};
  assign memory[349] = {`SW, `SP, `A1, 16'd16};
  assign memory[350] = {`SW, `SP, `A2,  16'd20};
  assign memory[351] = {`SW, `SP, `RA,  16'd24};
  assign memory[352] = {`NOP};
  assign memory[353] = {`ADDI, `ZERO, `T1, 16'd0}; //T1 is the loop counter
  assign memory[354] = {`ADDI, `ZERO, `T2, 16'd6};
  assign memory[355] = {`J, 26'd376}; //condition
  assign memory[356] = {`NOP};
  assign memory[357] = {`NOP};
  assign memory[358] = {`NOP};
  assign memory[359] = {`NOP};
  assign memory[360] = {`NOP}; // for_body
  assign memory[361] = {`LW, `SP, `T4, 16'd0};		//x coordinate
  assign memory[362] = {`LW, `SP, `T5,  16'd4};		//y coordinate
  assign memory[363] = {`ADDI, `T5, `T6, 16'd1}; 	//increment y coordinate
  assign memory[364] = {`LW, `SP, `A0,  16'd8};		//color
  assign memory[365] = {`SPECIAL, `NULL, `A0, `A0, 5'd16, `SLL};
  assign memory[366] = {`ORI, `A0, `A0, `T4, `T5};
  assign memory[367] = {`JAL, 26'd418}; //write_byte
  assign memory[368] = {`ADDI, `T1, `T1, 16'd1}; //increment loop counter
  assign memory[369] = {`SW, `SP, `T6, 16'd4}; //update x coord. counter
  assign memory[370] = {`NOP};
  assign memory[371] = {`NOP};
  assign memory[372] = {`NOP};
  assign memory[373] = {`NOP};
  assign memory[374] = {`NOP};
  assign memory[375] = {`NOP};
  assign memory[376] = {`NOP}; //condition
  assign memory[377] = {`SPECIAL, `T1, `T2, `T3, `NULL, `SLT};
  assign memory[378] = {`BNE, `T3, `ZERO, 16'ha}; // for_body
  assign memory[379] = {`NOP};
  assign memory[380] = {`LW,`SP,`A0,  16'd12};
  assign memory[381] = {`LW,`SP, `A1,  16'd16};
  assign memory[382] = {`LW,`SP, `A2,  16'd20};
  assign memory[383] = {`LW,`SP, `RA, 16'd24};
  assign memory[384] = {`NOP};
  assign memory[385] = {`ADDI, `SP, `SP, 16'd32};
  assign memory[386] = {`SPECIAL, `RA, 15'd0, `JR};
  assign memory[387] = {`NOP};
  assign memory[388] = {`NOP};
  assign memory[389] = {`NOP};
  assign memory[390] = {`NOP}; //pause
  assign memory[391] = {`ADDI, `ZERO, `T0, 16'd0};
  assign memory[392] = {`ADDI, `ZERO, `T1, 16'h100};
  assign memory[393] = {`J, 26'd412}; //pause_outer_condition
  assign memory[394] = {`NOP};
  assign memory[395] = {`NOP};
  assign memory[396] = {`NOP}; //pause_outer
  assign memory[397] = {`ADDI, `T0, `T0, 16'd1};
  assign memory[398] = {`ADDI, `ZERO, `T4, 16'd0};
  assign memory[399] = {`ADDI, `ZERO, `T5, 16'd1};
  assign memory[400] = {`J, 26'd407}; //pause_inner_condition
  assign memory[401] = {`NOP};
  assign memory[402] = {`NOP};
  assign memory[403] = {`NOP}; //pause_inner
  assign memory[404] = {`ADDI, `T4, `T4, 16'd1};
  assign memory[405] = {`NOP};
  assign memory[406] = {`NOP};
  assign memory[407] = {`NOP}; //pause_inner_condition
  assign memory[408] = {`SPECIAL, `T4, `T5, `T6, `NULL, `SLT};
  assign memory[409] = {`BNE, `T6, `ZERO, 16'ha}; //pause_inner
  assign memory[410] = {`NOP};
  assign memory[411] = {`NOP};
  assign memory[412] = {`NOP}; //pause_outer_condition
  assign memory[413] = {`SPECIAL, `T0, `T1, `T2, `NULL, `SLT};
  assign memory[414] = {`BNE, `T2, `ZERO, 16'ha}; //pause_outer
  assign memory[415] = {`SPECIAL, `RA, 15'd0, `JR};
  assign memory[416] = {`NOP};
  assign memory[417] = {`NOP};
  assign memory[418] = {`NOP}; //function: write_byte
  assign memory[419] = {`ADDI, `ZERO, `T0, 16'hffff};
  assign memory[420] = {`SPECIAL, `NULL, `T0, `T0, 5'd16, `SLL};
  assign memory[421] = {`SW, `T0, `A0, 16'hc};
  assign memory[422] = {`SPECIAL, `RA, 15'd0, `JR};
  assign memory[423] = {`NOP};
  assign memory[424] = {`NOP};
  assign memory[425] = {`NOP};
  assign memory[426] = {`NOP};
  assign memory[427] = {`NOP};
  assign memory[428] = {`NOP};
  assign memory[429] = {`NOP};
  assign memory[430] = {`NOP}; // poll_for_ready
  assign memory[431] = {`LW, `T8,`T9,  16'd20};
  assign memory[432] = {`ANDI ,`T9, `T9, 16'd1};
  assign memory[433] = {`BLEZ, `T9, 5'b0, -16'd4}; //poll_for_ready 
  assign memory[434] = {`NOP};
  assign memory[435] = {`SW, `T8, `A0,  16'd4};
  assign memory[436] = {`SPECIAL, `RA, 15'd0, `JR};
  assign memory[437] = {`NOP};
  assign memory[438] = {`NOP};
  assign memory[439] = {`NOP}; //end_the_game
  assign memory[440] = {`ADDI, `ZERO, `A0, 16'd69}; // 69 is 'E'
  assign memory[441] = {`JAL, 26'd418}; //jump to write_byte
  assign memory[442] = {`NOP};
  assign memory[443] = {`ADDI, `ZERO, `V0, 16'd10}; //the exit syscall
  assign memory[444] = {`NOP}; 
  assign memory[445] = {`NOP};
  assign memory[446] = {`NOP};
  assign memory[447] = {`NOP};
  assign memory[448] = {`NOP};
  assign memory[449] = {`NOP};
  assign memory[450] = {`NOP};
  assign memory[451] = {`NOP};
  assign memory[452] = {`NOP};
  assign memory[453] = {`NOP};
  assign memory[454] = {`NOP};
  assign memory[455] = {`NOP};
  assign memory[456] = {`NOP};
  assign memory[457] = {`NOP};
  assign memory[458] = {`NOP};
  assign memory[459] = {`NOP};
  assign memory[460] = {`NOP};
  assign memory[461] = {`NOP};
  assign memory[462] = {`NOP};
  assign memory[463] = {`NOP};
  assign memory[464] = {`NOP};
  assign memory[465] = {`NOP};
  assign memory[466] = {`NOP};
  assign memory[467] = {`NOP};
  assign memory[468] = {`NOP};
  assign memory[469] = {`NOP};
  assign memory[470] = {`NOP};
  assign memory[471] = {`NOP};
  assign memory[472] = {`NOP};
  assign memory[473] = {`NOP};
  assign memory[474] = {`NOP};
  assign memory[475] = {`NOP};
  assign memory[476] = {`NOP};
  assign memory[477] = {`NOP};
  assign memory[478] = {`NOP};
  assign memory[479] = {`NOP};
  assign memory[480] = {`NOP};
  assign memory[481] = {`NOP};
  assign memory[482] = {`NOP};
  assign memory[483] = {`NOP};
  assign memory[484] = {`NOP};
  assign memory[485] = {`NOP};
  assign memory[486] = {`NOP};
  assign memory[487] = {`NOP};
  assign memory[488] = {`NOP};
  assign memory[489] = {`NOP};
  assign memory[490] = {`NOP};
  assign memory[491] = {`NOP};
  assign memory[492] = {`NOP};
  assign memory[493] = {`NOP};
  assign memory[494] = {`NOP};
  assign memory[495] = {`NOP};
  assign memory[496] = {`NOP};
  assign memory[497] = {`NOP};
  assign memory[498] = {`NOP};
  assign memory[499] = {`NOP};
  assign memory[500] = {`NOP};
  assign memory[501] = {`NOP};
  assign memory[502] = {`NOP};
  assign memory[503] = {`NOP};
  assign memory[504] = {`NOP};
  assign memory[505] = {`NOP};
  assign memory[506] = {`NOP};
  assign memory[507] = {`NOP};
  assign memory[508] = {`NOP};
  assign memory[509] = {`NOP};
  assign memory[510] = {`NOP};
  assign memory[511] = {`NOP};

endmodule
